--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:44:55 12/13/2013
-- Design Name:   
-- Module Name:   C:/hlocal/toc/Practica5/practica5/miTest.vhd
-- Project Name:  practica5
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: practica5
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY miTest IS
END miTest;
 
ARCHITECTURE behavior OF miTest IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT practica5
    PORT(
         rst : IN  std_logic;
         clk : IN  std_logic;
         inicio : IN  std_logic;
         fin : OUT  std_logic;
         direccion : IN  std_logic_vector(4 downto 0);
         dato_debug : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal rst : std_logic := '0';
   signal clk : std_logic := '0';
   signal inicio : std_logic := '0';
   signal direccion : std_logic_vector(4 downto 0) := (others => '0');

 	--Outputs
   signal fin : std_logic;
   signal dato_debug : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: practica5 PORT MAP (
          rst => rst,
          clk => clk,
          inicio => inicio,
          fin => fin,
          direccion => direccion,
          dato_debug => dato_debug
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      rst<='1';
      wait for 100 ns;	
		rst<='0';
		wait for clk_period;
		inicio <= '1';
      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
