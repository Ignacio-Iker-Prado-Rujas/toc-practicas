--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   19:16:20 11/29/2013
-- Design Name:   
-- Module Name:   C:/hlocal/toc-practicas/Practica4/prueba1.vhd
-- Project Name:  Practica4
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: maquina_divisor
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY prueba1 IS
END prueba1;
 
ARCHITECTURE behavior OF prueba1 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT maquina_divisor
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         divisor : IN  std_logic_vector(7 downto 0);
         dividendo : IN  std_logic_vector(15 downto 0);
         inicio : IN  std_logic;
         ready : OUT  std_logic;
         cociente : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal divisor : std_logic_vector(7 downto 0) := (others => '0');
   signal dividendo : std_logic_vector(15 downto 0) := (others => '0');
   signal inicio : std_logic := '0';

 	--Outputs
   signal ready : std_logic;
   signal cociente : std_logic_vector(15 downto 0);

   -- clk period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: maquina_divisor PORT MAP (
          clk => clk,
          reset => reset,
          divisor => divisor,
          dividendo => dividendo,
          inicio => inicio,
          ready => ready,
          cociente => cociente
        );

   -- clk process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		dividendo <= "1011010110101010";
		divisor <= "10101001";
		
      wait for clk_period*10;
		
		inicio <= '1';
		
		wait for 100 ns;

      -- insert stimulus here 

      wait;
   end process;

END;
